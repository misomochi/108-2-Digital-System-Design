`timescale 1ns/10ps
`define CYCLE  10
`define HCYCLE  5

module register_file_tb;
    // port declaration for design-under-test
    reg        Clk, WEN;
    reg  [2:0] RW, RX, RY;
    reg  [7:0] busW;
    wire [7:0] busX, busY;

    parameter count = 8;
    integer i, err;
    
    // instantiate the design-under-test
    register_file rf(
        Clk  ,
        WEN  ,
        RW   ,
        busW ,
        RX   ,
        RY   ,
        busX ,
        busY
    );

    // write your test pattern here
    initial begin
        $fsdbDumpfile("register_file.fsdb");
        $fsdbDumpvars;
    end

    always #(`HCYCLE) begin
        Clk = ~Clk;
    end

    initial begin
        Clk  = 0;
        WEN  = 0;
        RW 	 = 0;
        RX 	 = 0;
        RY 	 = 0;
        busW = 0;
        err = 0;

    	for (i = 0; i < count; i = i + 1) begin
    		@(negedge Clk);
    		WEN = 1;
    		RW = i;
    		busW = $unsigned($random) % 8'b1111_1111;
    		$display("Write %b to reg %d.", busW, RW);

    		@(negedge Clk);
    		WEN = 0;
    		RX = i;
    		RY = i;

    		@(negedge Clk);
    		if (i == 0) begin
    			if (busX !== 8'b0 || busY !== 8'b0) begin
    				$display("ERROR at reg %d: X output %b != %b", RX, busX, 8'b0);
    				$display("ERROR at reg %d: Y output %b != %b", RY, busY, 8'b0);
    				err = err + 1;
    			end
    			else begin
    				$display("%d-th test PASSED: X output %b == %b", RX, busX, 8'b0);
    				$display("%d-th test PASSED: Y output %b == %b", RY, busY, 8'b0);
    				err = err;
    			end
    		end
    		else begin
    			if (busX !== busW || busY !== busW) begin
    				$display("ERROR at reg %d: X output %b != %b", RX, busX, busW);
    				$display("ERROR at reg %d: Y output %b != %b", RY, busY, busW);
    				err = err + 1;
    			end
    			else begin
    				$display("%d-th test PASSED: X output %b == %b", RX, busX, busW);
    				$display("%d-th test PASSED: Y output %b == %b", RY, busY, busW);
    				err = err;
    			end
    		end
    	end

    	if (err == 0) begin
    		$display("                                                                                   *****************//&&&&&&@&#&/&(/*****************************/    ");
			$display("                                                                                   *********************#/&/..#&@/@*&,@/&&#/*/*******************/    ");
			$display("                                                                        ,,,*,,*****(*******,*********************(#//(..#&&&&&&#*****************(    ");
			$display("                                                                    ,,,,*,,,,,,,,,,,,**/*,*****************,,*,,,******///(/&&&//****************#    ");
			$display("        *******//*/*   /*/*,                                     ,*,,,,,,,,,,,,......,,*,**/*******,**********,,*,*,*,**************************/     ");
			$display("               *///    ////                                    *,,.......,,...........,,,,,,//************,***,,,*******************************      ");
			$display("         **    *///   */*/                                    *,,....................,,,,,,,*//,**********,**,,********/*******,***************       ");
			$display("         ////  ,//*   *//,                                   *,,,,,................,,,,,,,,,,*/,,*********,*,,*,,,***********************,***(        ");
			$display("         /*/.  .//.   */* /*                                .*,,,,,................,,,,,,,,,**//,********,,,,*,,,*,*******,*****************.         ");
			$display("         ///   **//  *//   ///                              ***,,,,......,.,,,,.,,,,,,,,,,,,**/(,,**(//(#/***//*(************************/&           ");
			$display("               /*/,  //     ///,                            /***,,,,,,,,.,,**,,,,,,****,,,,***/(,*#//*@@@@@&@*@#*/(//****,**********,*(&#             ");
			$display("               /*/  **,*////////                            //(((((((((*,,,,//((#/#((///,,,***/(.(,*@&@#@@@&&@/@/@*(*********,*****#&##               ");
			$display("           .*//*/.//*//,     //*                           .*/((**##,/*/,.,*,,.,,,.,,****,,**/(***,@&&&@#&/&&&&@@@@*((**********/#@                   ");
			$display("             ,.                                            ,//*,,,,,,,**,.,,*,......,,,,,,,**/*,,.*&&&&&&&&,&/&@&&@,#*,,******,(                      ");
			$display("                                                           .**,.....,*/,,.,,**,.......,,,******,**(*&#&&&&&&/&#&&&,#,***,*,***&                       ");
			$display("          *//*      *///,                                  ,/*,,,,,****,..,,*,/**,,,,,,**/*///,*,*//(//@(&@&&#&&*/(**,,*,,,,,,/                       ");
			$display("            **/.    */*/                                    (((////**(/////#(/*,,,*(/////*//((*,***/##*#///&&(#(*&,**,*,,,****/                       ");
			$display("               **//*//*/*///*/*                             /(/*,//(******,,,,,**/(/*,****/#(//***///#//#&,/#//*****,,,,******,.                      ");
			$display("         ///* /.    */*/                                     (//*,,,/*//*,******,...,****/(((*/*///////(#// (/**,***,***,*,,*,,/                      ");
			$display("          ,/ /,     ///*    /*,                                (/((**,***/**,,,.,,*/**/(#/******/*(//#**///&/*********,*,*,***,/                      ");
			$display("           ./*     /*///                                         /##/***,..,,****(#((#/&***,*****#/##*#/*///***,*,**********,,*                       ");
			$display("          ///     ///*  /*                                         /&/(((//((/(#&//&&/**,,,****/,//**///&*//**,***,**,********                        ");
			$display("          */*    **,      ///,                                     ***/###//&&&/(///**,,,,****/**.(/&/&////*********,******(*                         ");
			$display("          ////***/////*    ///*                                 ,#*****(///,,,.,,,,,,,,,,****/**///&/&//////*/*********/#&                            ");
			$display("           *,  *.           *.                             ,**,#/(******(//*,,,,,,,,.,,,******,&//////#*,,,,#&&&&&&&&(*                               ");
			$display("                                                      .*,,,,,*#/***********//**,,,,.,,***,*,,,/&//&*(///,,,,,,,,,,,,,,,,***.                          ");
			$display("                                                   .,,,*,,,,(#*,************,,,,,,,..***,,,,,##,(/&&#/&,,,,,,,,,,,,,,,,,,,,,*,.                       ");
			$display("              //*     ///   //                   ,,,***,**,##**,,********,**,..,,,,.*,,,,,,,,(//**/#//(,,,,,,,,,,,,,,,,,,,,,,,,*.                     ");
			$display("              //*     //*                       ,,,/*,,,,,//*,,,,,,,**,,,*,,,*,,,,,,,,,,,,,,/&//&(//,(/,,,,,,,,,,,*,,,**,,,,,,,,**                    ");
			$display("              //*     //,                     ,,*,/*,,,,/#/*,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,/.*//&&/&/#*,,,,,,,,,,,*,,**,,,,,,,,,,,,*                  ");
			$display("              */,    *//*/                   ***,*,,,,,/*(*,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,(/////,//((*,,,,,,,,,,,*,,*,,,,,,,,,,,,*,,                 ");
			$display("           ///, */  .///.                   .*,,,,,,,,*/#*,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,/&//,/&&#(#/*,,,,,,,,,,**,**,,,,,,,,,,,,*,*,                ");
			$display("           //    /*//**                     **,,,,,,,,##*,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,//&/(&&//##,*,,,,,,,,,,**,/,,,,,,,,,,,,,,,,,,               ");
			$display("                 *///*/                    .*,*,,*,,,(/**,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,#&&(//.#/,#(,*,,,,,,,,,,*,,*,,,,,,,,,,,,*,,,,,,              ");
			$display("              ,//*,  ///*///*,.            ***,,,,,,*//*,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,/&///#&&&,*//,*,,,,,,,,,****,,,,,,,,,,,,,,,,,*,*.             ");
			$display("          .///.         ,/////             **,,*,,,*#(*,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,/&&/#&#,,**/*,,*,,,,,,,,***,,,,,,,,,,,,,*,,,,*,,/             ");
			$display("                                          .********/#**,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,#&&#/&/&/,/*((,,*,,,,,,,,**,,,,,,,,,,,,,*,,,,,*,,,/            ");
			$display("                                          **********,**,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,/&#&&#/*/,/(#,/,,,,,,,,,,,**,*,,,,,,,,,,,*,,,***,*,*/           ");
			$display("          ///*       //*/   .             ********/(**,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,#&&&#&&/,,((**//,,,,,,,,*,*,*,*,,,,,,,,***,****,*****,          ");
			$display("         //** .******///*******          ***/****##((**,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,/&&#&#,(/,#/(,,/(**,,,,********,,,*********,*********,*          ");
			$display("        *. ,,  ***///////////*,          (*//*/*(###/**,,,,,,,,,,,,,,,,,,,,,,,,,,,,,/&#&&&(&&,*/(,**/##*,,,*****,*,*,**/********,***,*,*,****         ");
			$display("          *///.*//,,// //* ///          ,/***////###***,****,,,,,,,,,,,,,,,,,,,,,,,,#&&,*&&(,,(*(,,/#*/*,,******,*****/********************/*,        ");
			$display("         ////  **/**//*///*/*/          ///*///#/###********,,,,,,,,,,,,,,,,,,,*,,,&&&#&&&(,,*##*,*/#*(*********,****/******************,,/***        ");
			$display("        ////,              ,//*        ,*//*(*/#*(#/********,*,,,,,,,,,,,,,,,,,,,,,/#&&&*&/,,#/#,**((*##************/********************/*****       ");
			$display("         ///.        //*               /*****/(#(*(/********,,,,,,,,*,,,,,,,,,,*,//&&&#&  ,,*##**,#(#(##(*****/****/******************,********       ");
			$display("         ///. */ */** .// / ///       ./*****(/(#**#/*******,,,,,,,,*,,*,,,,,,,(&/,/&&/./&,,#(/*,*####(##****//***//**********************///(*,      ");
			$display("         ///./// *///*////* ./*       //*****###(**#/********,,*,****,,,,,,,,/(&.*/&&&*,*&*#(/*,**#######***///**///****(/*************//((/***,      ");
			$display("         /*/      .*******,           //****/##(***#/*********,*,****,,,,,,**,&/,,#&&, .&/&//****(#####/#****///*(//**/(*************/#/********      ");
			$display("                                     ,//****/((#***#(********,,***,**,,,,,,*/&//*,&&&***&*##(*,*,#/####/#*****///(/****//(#((((/***/**********/,      ");
			$display("                                     ,/(/***((#/***##*/**************,,***,,/&,**&&&..,&##//***,/###(#////*/**************,**,****/**********//.      ");
			$display("                                     ./(/***###****(#*/*************,*,,,,//&***#(********,,,,,*,*,,,,,*,,,,,***,,/**************************/(.      ");
			$display("                                      ((/***##(****(#(/*,,,*,,,...,,,,,,*,,,,,,,,,,,,,,,,,*/,,***,,,,,,,**,*,,,*,,***************************/(       ");
			$display("                                      ((/*/(##*****/(#/**#(/*//*,....,,,,,,,,,,,,,,,,,,,,,,******,,,,*,**,********,***************//*/////////(       ");
			$display("                                      ,(/**##(*****/(#/***/,,,***,...,,******************************************/**********///////////////////       ");
    	end
    	else begin
    		$display(" .,,**,,,,*//**********,....                            ..    .....,,,,*****////((((((((((((#(#####(");
			$display(" ....,**,,,,,***,,..                                  .     .............,,*//((((/((#//#/****/(#(/*");
			$display(" .,***/*,,,,,..                           .       .........................,,*////////((////****////");
			$display(" ......,,...                    ..   ......     ............................,,,,,**///////*//(/*////");
			$display("  ............          /@@@@@@@& @@@@@@@@ @@@@.@@@@..@@@@@@@@.@@@@..@@@@@@@@ ,,,,,,****************");
			$display("  ....   .....          @@@@ @@@@...@@@@...@@@@.@@@@,.@@@, @@@,@@@@..@@@* @@@&,,,,,,,*/(((/*//*,,***");
			$display("......   ................@@@@@@.....@@@@...@@@@.@@@@,.@@@@@@@@,@@@@, @@@* @@@@,,,.....,,,,****,,,,,*");
			$display(".....    ...............    *@@@@.. @@@@...@@@@.@@@@..@@@, ....@@@@..@@@* @@@@..........,******,,,,,");
			$display("...      ...............@@@@.@@@@   @@@@.. @@@@ @@@@..@@@,     @@@@. @@@*.@@@/ ** ........,*//****,,");
			$display("           ...       ... *@@@@@@   .@@@@    #@@@@@&  .@@@,     @@@@  @@@@@@@/  @@... ......*(/**//**");
			$display("                                                                            .  ....     .. .,*//////");
			$display("                                                                                         ....,**/**/");
			$display("                                                                                        .....,*/(###");
			$display("                                                  ..   ..                      ..    ... ..  .,*****");
			$display("                                             .............   .        ..   ..............    .,*****");
			$display("                                  .....................,.........     ....................    .*////");
			$display("                                .....,,,,........,,,.,,,,,..................,,,,,,,........   .,////");
			$display("                                ..,,,,,,,,,,...,,,,,,,**,,,,...........,,,,,*********,,,,,,.  .,*///");
			$display("                              ....,,,********,,,,,***********,**********************//**///,  .,*///");
			$display("                          .......,,,,*******************////////////////////////////////(((*. .*///(");
			$display("                         .....,,,,************/////////////////////////////////////////////*,,,*****");
			$display("                        ....,,,*************/////////*/****///////////////************,,...,,***///*");
			$display("                        ....,,***********/////////****,,,......,,,*****************,,....,,***//////");
			$display("                        ...,,********/////////****,,,,,,,,,..........,**********,,,,,,,,****//##(///");
			$display("                       ....,*******////////************//****,,,,,,,,,,,*******,,,,,,,,......*((/*//");
			$display("                     .....,,,***//////////********,,,,.........,,,,,,,,*********,,,..   .,**,*((////");
			$display("           ...............,,,***//////////****,,,...,..   .,*,,..,,,******//****,,,,,,,,*****/(((((#");
			$display("  .,*/(///(/**,,..........,,****//////////*************,,****,,,,,******/////*****,,,,,,,*****/(/*//");
			$display(" .*/*,,.,,,,*****,,,......,,***//////////////////*********,,,,,,******//////////******,,,,****/(////");
			$display(",***,,*****,,,**,,,,,,...,,,*****/////////////////*********,,,******///////////(/************///////");
			$display("*///***//////**,,,,,**,,.,,,,*******////////////////***********//**********///((((/*******//////////");
			$display(",///////(//*,..,,,,*****,,,,,,,*******////////////////******/////**********////(((((/*****//////////");
			$display(".,*////(//*,,,,,,,,*//***,,,,,,**********/*****////////////////***********/////////(//****//////////");
			$display(" .,///////******,,,,******,,,,,,,,*********************/////**********///////*******///*******//((((");
			$display("  .*/(((////*******,,,******,,,,,,,,,,,,,,**************//*************/***,,,,,,,,,,,**************");
			$display("  .,/((/////////((//********,,,,,,,,,,,,,,,,,,********************,,,,,,............,,**********//**");
			$display("  .,//**/////((((//////*,,***,,,,,,,,,,,,,,,,,,,***************//***,.....,,,,,,,,,*****************");
			$display("  .,*/*,,,**//(((((((///*****,,,*,,,,,,,,,,,,,,,,,************/////***/**************/*******/(#//#(");
			$display("  .,/(((/,.....,*////////**,,,,,,,,,,,,,,,,,,,,,,,,*********************////*******************(#/**");
			$display("   .,,,,....      ...,,,....,,,****,,,,,,,,,,,,,,,,,,*********************,,,,,,,,....,,,******(#/**");
			$display("   .........       ..,,,,,...,,,*,*,,,,,,,,,,,,,,,,,,,********,,,,,,,,,......,,,......,,***////(#(//");
			$display("            .       .,,,,,,,..,,,,,,,,,,,,,,,,,,,,,,,,,***,,,,,,.        ..........,,*,*****///***//");
			$display("            ...     ..,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,*,,,,,,,,,,,,,,,,,,,,,******************//");
			$display("               ....  ...,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,,***,,,,,,,,,,,,,,*******************");
			$display("                .........,,,,,,,,,...,,,,,,,,,,,,,,,,,,,,,,,,,,,*,,,,,,,...,,,,,,,,****(#/#((#((###(");
			$display("                    ......,,,,,,,,.......,,,,,,,,,,,,,,,,,,,,*******,,,,........,,*************/##/*");
			$display("                      ......,,,,,,,...........,,,,,,,,,,,********************,*****************/##/*");
			$display("                         .....,,,,,..............,,,,,,,*********************************///////##(/");
			$display("                           ......,....................,,,,,**************************//(/#(/////////");
			$display("                 .              .........................,,,,,,,,*********,,,,,,,,,,***/##/*********");
    	end

    	$finish;
    end

endmodule
